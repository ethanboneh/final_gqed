
// ------------------------------------------------------------------
//   Design Unit:    GQED_rtl
// ------------------------------------------------------------------


// We will check FC of read action
// Though there exists a solution such that the code apart from /*Fill*/ and /*Code goes here*/ needs no modification, feel free to modify the code as per convenience.

module gqed
#(
parameter SEQ_LEN = 32, // Maximum length of the pre-sequence. Pre-sequence is fed to both first and second copy.
RESP_BOUND = 2 // Upper bound estimate of the number of clock cycles for read action to finish execution 
)
(
// BMC controlled inputs

input clk, clk_en, rst,
input [$clog2(SEQ_LEN)-1:0] i, // index of input under verification in first copy. By definition, i<SEQ_LEN.
input [32:0] in [0:SEQ_LEN-1], // stores the pre-sequence and the input under verification [in[0],...in[i]]. First 16 bits (in[*][15:0]) is address, next 16 bits (in[*][31:16]) is data and the MSB (in[*][32]) decides action (read (in[*][32]==1'b0), write (in[*][32]==1'b1)).
input in_vld2, // BMC chooses input to be valid or invalid in the second copy. Note that BMC should be able to exercise all possible input sequences in the second copy. Otherwise, there will be completeness issues.
input [33:0] bmc_in2 // BMC gets to choose this input. Used in second copy when in_vld2 is low and for the inputs after in_i. bmc_in2[33:32] feeds ren_in and wen_in separately. 
);

reg [7:0] bound; // Wait for RESP_BOUND clock cycles after i-1 inputs have been fed to first copy.  
 
reg [$clog2(SEQ_LEN)-1:0] cntr1, cntr2, cntr3; // keeps track of sequence index of the inputs being fed to the three copies. 
reg [$clog2(SEQ_LEN)-1:0] ocntr2; // keeps track of the sequence index of the outputs generated by the second copy. Output is only generated by read actions.
reg [$clog2(SEQ_LEN)-1:0] no_ocntr2; // keeps track of the number of inputs that produce no output i.e. inputs with write action (in[*][32]==1'b1).  


reg [15:0] arch_st1_i; // saves value of the arch state after idling in the first copy.
reg [15:0] arch_st3_i; // saves value of the arch state right after reset in the third copy. 

reg arch_st_done1, arch_st_done3; // goes high when the arch state is saved in first and third copies.

reg [15:0] cmp_out2, cmp_out3; // out2 saves i^th output from the second copy, out3 saves 1st output in the third copy. The first input in the third copy is the same as the i^th input in the second copy. 

reg done2, done3; // goes high when output is saved in second and third copies.

reg ren_d2, ren_d3; // signals to look at the value of the ren_in signal one clock cycle before for the second and third copies. The output is generated after 1 clock cycle since the read action is fed. 


//ports to interface with the three copies
wire [15:0] addr_in1, data_in1, addr_in2, data_in2, out2, addr_in3, data_in3, out3; 
wire wen_in1, ren_in1, wen_in2, ren_in2, wen_in3, ren_in3; 


//instantiation of the 3 copies
memory_core copy1 (.clk(clk), .clk_en(1'b1), .reset(rst), .flush(1'b0), .config_en_sram(4'b0), .enable_chain(1'b0), .tile_en(1'b1), .addr_in(addr_in1), .data_in(data_in1), .wen_in(wen_in1), .ren_in(ren_in1), .mode(2'd2));
memory_core copy2 (.clk(clk), .clk_en(clk_en), .reset(rst), .flush(1'b0), .config_en_sram(4'b0), .enable_chain(1'b0), .tile_en(1'b1), .addr_in(addr_in2), .data_in(data_in2), .wen_in(wen_in2), .ren_in(ren_in2), .mode(2'd2), .data_out(out2));
memory_core copy3 (.clk(clk), .clk_en(1'b1), .reset(rst), .flush(1'b0), .config_en_sram(4'b0), .enable_chain(1'b0), .tile_en(1'b1), .addr_in(addr_in3), .data_in(data_in3), .wen_in(wen_in3), .ren_in(ren_in3), .mode(2'd2), .data_out(out3));


assume property (@(posedge clk) in[i][32] == 1'b0); // we will check FC of read action only. 


  /*
     Write constraints for input signals and the arch state. in and i needs to be held constant. The arch state right after reset should be the same for the first and second copies otherwise even the same input preseqeuence will not guarantee same arch state.
     Signals to use: i, in, rst,  copy1.mem_inst0.sram_stub.data_array, copy1.mem_inst1.sram_stub.data_array, copy2.mem_inst0.sram_stub.data_array, copy2.mem_inst1.sram_stub.data_array
  */  

stable_in: assume property (@(posedge clk) $stable(in));
stable_i: assume property (@(posedge clk) $stable(i));
same_arch_state_at_rst: assume property (@(posedge clk) $fell(rst) |-> copy1.mem_inst0.sram_stub.data_array == copy2.mem_inst0.sram_stub.data_array && copy1.mem_inst1.sram_stub.data_array == copy2.mem_inst1.sram_stub.data_array);

// ------------------------------------------------------------------   


  /*
     Write constraints for input signals and the arch state. in and i needs to be held constant. The arch state right after reset should be the same for the first and second copies otherwise even the same input preseqeuence will not guarantee same arch state.
     Signals to use: i, in, cntr1, in_vld2, cntr2, bmc_in2
  */ 

// copy 1

assign addr_in1 = in[cntr1][15:0]; // read data from in based of counter position. 
assign data_in1 = in[cntr1][31:16]; // similarly read address 

  /*
     To write, wen_in has to be high. We don't care about ren_in (1'bx). To read, wen_in == 1'b0 and ren_in == 1'b1. After i-1 inputs, we have to idle i.e. no valid inputs (wen_in == 1'b0 and ren_in == 1'b0). 
     Hint: can use nested ternary operators 
  */

assign wen_in1 =  cntr1<i? in[cntr1][32]:1'b0; 
assign ren_in1 = cntr1<i?(in[cntr1][32]?1'bx:1'b1):1'b0; 
// ------------------------------------------------------------------   

// copy 2

  /*
     Fill in similar to first copy. Now we have to send the first i inputs from in. If BMC decides to send an invalid input (in_vld2 == 1'b0) and for inputs after i^th input, feed from bmc_in2. 
  */

assign addr_in2 = in_vld2 && cntr2<=i?in[cntr2][15:0]:bmc_in2[15:0];
assign data_in2 = in_vld2 && cntr2<=i?in[cntr2][31:16]:bmc_in2[31:16];
assign wen_in2 = in_vld2 && cntr2 <= i? in[cntr2][32] : (cntr2 <= i ? 1'b0 : bmc_in2[33]);
assign ren_in2 = in_vld2 && cntr2 <= i? (in[cntr2][32]?1'bx:1'b1) : (cntr2 <= i ? 1'b0 : bmc_in2[32]);
// ------------------------------------------------------------------   

// copy 3

  /*
     Fill in similar to first copy. We only care about the first input, the j^th input from in. 
  */

assign addr_in3 = in[i][15:0];
assign data_in3 = in[i][31:16];
assign wen_in3 = cntr3<1?in[i][32]:1'b0;
assign ren_in3 = cntr3<1?(in[i][32]?1'bx:1'b1):1'b0;

// ------------------------------------------------------------------   


  /*
     Logic for input index tracking counter in the second copy. If the input is valid, increment cntr2. Update no_ocntr2 if the valid input is a write action. Make sure to prevent the counters from overflowing. 
     Signals to use: clk_en, in_vld2, cntr2, i, in    
  */

always @(posedge clk) begin
	if(rst) begin
		cntr2 <= 'b0;
		no_ocntr2 <= 'b0;
	end else begin 
		if (clk_en && in_vld2 && cntr2<=i) begin
			cntr2 <= cntr2 + 'b1;
			if (in[cntr2][32])
				no_ocntr2 <= no_ocntr2 + 'b1;
		end 			
	end
end

// ------------------------------------------------------------------   

  /*
     Logic for input index tracking counter in the first and third copies. Invalid inputs are fed in the first copy right after i-1 inputs are sent and in the third copy after 1st input is sent. We also need to save arch state after the waiting for RESP_BOUND clock cycles after i-1 inputs are sent in the first copy and right after reset in the third copy. Note that clock is always enabled in the first and third copies. Make sure to prevent the counters from overflowing. Note that the MSB of the address is used to select between mem_inst0 (MSB == 0) and mem_inst1 (MSB == 1) and remaining 8 bits to map to access elements in the mem_inst0.sram_stub.data_array (size 512 elements each element 16 bits long).   
     Signals to use: cntr1, i, bound,  copy1.mem_inst1.sram_stub.data_array, copy1.mem_inst0.sram_stub.data_array, copy2.mem_inst1.sram_stub.data_array, copy2.mem_inst0.sram_stub.data_array      
  */

always @(posedge clk) begin
	if(rst) begin
		cntr1 <= 'b0;
		cntr3 <= 'b0;
		bound <= 'b0;
		arch_st_done3 <= 1'b0;
		arch_st_done1 <= 1'b0;
	end else begin 
		if (cntr1<i)
			cntr1 <= cntr1 + 'b1;
		if (cntr1 == i && bound < RESP_BOUND-1 && i>0)
			bound <= bound + 'b1;			
		if (bound == (i==0?0:RESP_BOUND-1)) begin
			if(in[i][9])
				arch_st1_i <= copy1.mem_inst1.sram_stub.data_array[in[i][8:0]];
			else
				arch_st1_i <= copy1.mem_inst0.sram_stub.data_array[in[i][8:0]];
			arch_st_done1 <= 1'b1;									
		end 

		if (cntr3<1) begin
			cntr3 <= cntr3 + 'b1;
			if(cntr3==0) begin
				if(in[i][9])
					arch_st3_i <= copy3.mem_inst1.sram_stub.data_array[in[i][8:0]];
				else
					arch_st3_i <= copy3.mem_inst0.sram_stub.data_array[in[i][8:0]];
				arch_st_done3 <= 1'b1;
			end						
		end 			
	end
end

// ------------------------------------------------------------------   


  /*
     Create logic for ren_d2 and ren_d3. Note that clk_en is always high in third copy. Remember that if wen_in is high, irrepsective of ren_in, the action will always be write so be sure to exclude that condition while updating ren_d*. ren_d* keeps track if the input in the last clock cycle was a valid read action or not. 
     Signals to use: in_vld2, in, cntr2, ren_in3      
  */

always @(posedge clk) begin
	if(rst)
		ren_d2 <= 1'b0;
	else if (clk_en)
		ren_d2 <= in_vld2 && !in[cntr2][32]; 
end

always @(posedge clk) begin
	if(rst)
		ren_d3 <= 1'b0;
	else 
		ren_d3 <= ren_in3; 
end

// ------------------------------------------------------------------   

  /*
     Create logic for incrementing ocntr2 and saving the i^th output in the second copy. The valid output for a read action action is produced 1 clock cycle later. ren_d2 captures this. Write action does not produce any output but all inputs upto i can have both write (captured in no_ocntr2) and read (i-no_ocntr2) actions so be sure to take that into account.  
     Important signals to use: clk_en, ren_d2, ocntr2, i, no_ocntr2     
  */

always @(posedge clk) begin
	if(rst) begin
		ocntr2 <= 'b0;
		done2 <= 1'b0;
	end else begin 
		if (clk_en && ren_d2 && ocntr2<=i)
			ocntr2 <= ocntr2 + 'b1;
		if (clk_en && ren_d2 && (ocntr2 == i - no_ocntr2) && !done2) begin
			cmp_out2 <= out2;
			done2 <= 1'b1;
		end
	end
end

// ------------------------------------------------------------------   

  /*
     Similarly Create logic for saving the 1st output in the third copy. 
     Important signals to use: cntr3, ren_d3, done3      
  */

always @(posedge clk) begin
	if(rst) begin
		done3 <= 1'b0;
	end else if (cntr3>=1 && ren_d3 && !done3) begin
		cmp_out3 <= out3;
		done3 <= 1'b1;
	end 
end
// ------------------------------------------------------------------   

  /*
     If arch states of first and third copies have been saved, constrain them to be equal. 
     Important signals to use: arch_st_done1, arch_st_done3, arch_st1_i, arch_st3_i   
  */

constraint_arch_state: assume property (@(posedge clk) arch_st_done1 && arch_st_done3 |-> arch_st1_i==arch_st3_i);

// ------------------------------------------------------------------   

  /*
     Check if i^th output from the second copy, 1st output from the third copy and the arch state in the first copy have been saved, the two outputs match. 
     Important signals to use: done3, done2, arch_st_done1, cmp_out3, cmp_out2     
  */

functional_consistency_check: assert property (@(posedge clk) done3 && done2 && arch_st_done1 |-> cmp_out3 == cmp_out2);


endmodule 
