

// have a RAM that is a 2D array storing X,y. Send X,y through valid controlled by formal tool
/*
another RAM stores read_values. 
*/